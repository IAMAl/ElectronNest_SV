///////////////////////////////////////////////////////////////////////////////////////////////////
//
//	ElectronNest
//	Copyright (C) 2024  Shigeyuki TAKANO
//
//  GNU AFFERO GENERAL PUBLIC LICENSE
//	version 3.0
//
//	Address Generation Unit for Global Buffer Memory
//	Module Name:	BRAM_AGU
//	Function:
//					Address Generation
//					supprt Strided Address and Base Address
//					Address is continuously generated by Affine Equation;
//						- Addr = Addr +/ Stride
//						- Initial Addr value is set by Base address
//						- Repeating until counter achieves to zero
//
///////////////////////////////////////////////////////////////////////////////////////////////////

module BRAM_AGU
	import pkg_bram_if::*;
#(
	parameter int WIDTH_ADDR   		= 14,
	parameter int WIDTH_LENGTH 		= 14,
	parameter int WIDTH_STRIDE 		= 14,
	parameter int WIDTH_BASE   		= 14
)(
	input							clock,
	input							reset,
	input							I_En,				//Flag: Enable to Work
	input							I_Set,				//Flag: Set Config
	input	[WIDTH_LENGTH-1:0]		I_Length,			//Vector Access-Length
	input	[WIDTH_STRIDE-1:0]		I_Stride,			//Stride Factor
	input	[WIDTH_ADDR-1:0]		I_Base,				//Base Address
	output	[WIDTH_ADDR-1:0]		O_Addr,				//BRAM Address
	output							O_Term				//Flag: Termination
);


	//// Configuration Registers									////
	logic	[WIDTH_LENGTH:0]		R_Length;
	logic	[WIDTH_STRIDE:0]		R_Stride;
	logic	[WIDTH_ADDR-1:0]		R_Addr;


	//// Output														////
	//	 Address
	assign O_Addr			= R_Addr;

	//	 Flag: Terminal
	assign O_Term			= I_En & ( R_Length == 1 );


	//// Vector Access Count										////
	//	 Actual Access-Length = I_Length + 1
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_Length		<= '0;
		end
		else if ( I_Set ) begin
			//Set Access Length
			R_Length		<= I_Length + 1'b1;
		end
		else if ( I_En ) begin
			//Count
			R_Length		<= R_Length - 1'b1;
		end
	end


	//// Setting Stride Factor										////
	//	 Actual Stride Factor = I_Stride + 1
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_Stride		<= '0;
		end
		else if ( I_Set ) begin
			//Set Stride Factor
			R_Stride		<= I_Stride + 1'b1;
		end
	end


	//// Access Address												////
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_Addr			<= '0;
		end
		else if ( I_Set ) begin
			//Set Base Address
			R_Addr			<= I_Base;
		end
		else if ( I_En ) begin
			//Increment by Stride
			R_Addr			<= R_Addr + R_Stride;
		end
	end

endmodule