///////////////////////////////////////////////////////////////////////////////////////////////////
//
//	ElectronNest
//	Copyright (C) 2024  Shigeyuki TAKANO
//
//  GNU AFFERO GENERAL PUBLIC LICENSE
//	version 3.0
//
//	Address Generation Unit
//		Module Name:	AddrGenUnit_Ld
//		Function:
//						Generate Series of Addresses used for Loading.
//						Before starting, the unit is set by configuration data.
//						The data are after attribute word of the config block.
//						Address is continuously generated by affine equation;
//							Addr = Addr +/- Stride
//							Initial Address is set by Base Address,
//							Repeat time is defined by Access Length
//						The unit has two contexts.
//							Primary context is used for one request coming from outer
//							Secondary context is used for loading in primary context
//							This function is used in external memory access
//
///////////////////////////////////////////////////////////////////////////////////////////////////

module AddrGenUnit_Ld
#(
	parameter int WIDTH_ADDR		= 8,
	parameter int WIDTH_LENGTH		= 8
)(
	input							clock,
	input							reset,
	input							I_Cond,				//Flag: Condition
	input							I_Set_Config,		//Setting Config
	input							I_Write_Switch,		//Switch for Writing
	input							I_Read_Switch,		//End of Loading then Switch
	input							I_En_AddrGen,		//Enable to Calc
	input							I_Decrement,		//Flag: Decriment for Address
	input	[WIDTH_LENGTH-1:0]		I_Length,			//Access Length
	input	[WIDTH_ADDR-1:0]		I_Stride,			//Stride Factor
	input	[WIDTH_ADDR-1:0]		I_Base,				//Base Address
	output	[WIDTH_ADDR-1:0]		O_Address,			//Address
	output	logic					O_RNo,				//Read-Context No.
	output	logic					O_Term				//Flag: End of Calc
);


	//// Logic Connect												////
	logic						EnUpdate;				//Enable Update
	logic [WIDTH_ADDR/2:0]		Stride;					//Stride Factor


	//// Capture Signal												////
	logic [WIDTH_LENGTH:0]		R_AccCount	[1:0];      //Access Counter
	logic [WIDTH_ADDR:0]		R_Stride	[1:0]; 		//Stride Factor
	logic [WIDTH_ADDR-1:0]		R_Address	[1:0]; 		//Address


	//// Context Number												////
	logic						R_WNo;
	logic						R_RNo;


	//// Context-Switch Timing										////
	//	 Read -witch is same or later timing of Write-Switch


	//// Enable Address Calc										////
	//	 I_R_Context_Switch can be high when it is note yet terminated
	//	 Updating address is used after the switch
	//	 This is happen in External RAM
	assign EnUpdate			= I_En_AddrGen & ( R_AccCount[ R_RNo ] != '0 );


	//// Select Stride Factor or Branch Distance					////
	//	 Most-Significant Half Word:	Branch Taken
	//	 Least-Significant Half Word:	Branch NOT Taken
	assign Stride			= ( I_Cond & I_Set_Config ) ?		I_Stride[WIDTH_ADDR-1:WIDTH_ADDR/2] :
								( ~I_Cond & I_Set_Config ) ?	'0 :
																'0;


	//// Memory Address												////
	assign O_Address		= R_Address[ R_RNo ];


	//// Termination												////
	assign O_Term			= ( R_AccCount[ R_RNo ] == 1 ) & I_En_AddrGen;


	////
	assign O_RNo			= R_RNo;


	//// Write Context Number										////
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_WNo			<= '0;
		end
		else if ( I_Write_Switch ) begin
			R_WNo			<= ~R_WNo;
		end
	end


	//// Read Context Number										////
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_RNo			<= '0;
		end
		else if ( I_Read_Switch ) begin
			R_RNo			<= ~R_RNo;
		end
	end


	//// Access Counter												////
	//	 Count the number of accesses
	//	 Generates O_Term flag when reachees zero
	always_ff @( posedge clock ) begin: ff_acccount
		if ( reset ) begin
			R_AccCount[0]	<= '0;
			R_AccCount[1]	<= '0;
		end
		else if ( I_Set_Config ) begin
			R_AccCount[ R_WNo ]	<= I_Length + 1'b1;
		end
		else if ( EnUpdate ) begin
			// Count by End
			R_AccCount[ R_RNo ]	<= R_AccCount[ R_RNo ] - 1'b1;
		end
	end


	//// Capture Stride Factor										////
	//	 Set "Value + 1, ex. "0" -> 1 this avoids a "while-loop"
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_Stride[0]	<= '0;
			R_Stride[1]	<= '0;
		end
		else if ( I_Set_Config ) begin
			R_Stride[ R_WNo ]	<= I_Stride[WIDTH_ADDR/2-1:0] + 1'b1;
		end
	end


	//// Access Address												////
	always_ff @( posedge clock ) begin
		if ( reset ) begin
			R_Address[0]	<= '0;
			R_Address[1]	<= '0;
		end
		else if ( I_Set_Config ) begin
			// Set Base Address
			R_Address[ R_WNo ]	<= I_Base;
		end
		else if ( EnUpdate & I_Decrement ) begin
			// Decriment by Stride
			R_Address[ R_RNo ]	<= R_Address[ R_RNo ] - R_Stride[ R_RNo ];
		end
		else if ( EnUpdate & ~I_Decrement ) begin
			// Increment by Stride
			R_Address[ R_RNo ]	<= R_Address[ R_RNo ] + R_Stride[ R_RNo ];
		end
	end

endmodule
